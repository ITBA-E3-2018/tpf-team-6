//This module will keep count seconds till it hits 60 or the rst signal is high
module seconds_counter(seconds,rst,clk);


